library ieee;
use ieee.std_logic_1164.all;

entity OOR is
	Port(		a_in, b_in : in std_logic_vector(7 downto 0);
				o : out std_logic_vector(7 downto 0));
end OOR;

architecture behavioral of OOR is
begin
	
	o <= a_in or b_in;

end behavioral;